module UART_TOP(
    input           clk,
    input           reset,
    input           f_write,
    input [7:0]     i_TxData,
    input           i_RxData,
    output          o_RxDone,
    output          o_TxD,
    output [7:0]    o_RxD
);

wire                        ;

UART_TX         Tx(
    .clk(clk),
    .reset(reset),
    .i_clk_tx(i_clk_tx),
    .i_switch(w_TxD),
    .TxStart(!empty),
    .TxDone(TxDone),
    .o_txd(o_TxD)
);

UART_RX         Rx(
    .clk(clk),
    .reset(reset),
    .i_clk_rx(i_clk_rx),
    .i_rxd(i_RxData),
    .RxDone(o_RxDone),
    .o_RxStopBit(),
    .o_rx_data(w_RxD)
);

FIFO            fifo(
    .clk(clk),
    .reset(reset),
    .rd(TxDone),
    .wr(f_write),
    .wr_data(wr_data),
    .empty(empty),
    .full(),
    .rd_data(rd_data)
);

clk_div         BRG(
    .clk(clk),
    .reset(reset),
    .o_clk_rx(o_clk_rx),
    .o_clk_tx(o_clk_tx)
);

endmodule